CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1358 699
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
76546066 0
0
6 Title:
5 Name:
0
0
0
28
13 Logic Switch~
5 50 443 0 1 11
0 22
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4484 0 0
2
5.90137e-315 0
0
13 Logic Switch~
5 49 420 0 1 11
0 24
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5996 0 0
2
5.90137e-315 0
0
13 Logic Switch~
5 51 390 0 1 11
0 25
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7804 0 0
2
5.90137e-315 0
0
13 Logic Switch~
5 52 361 0 1 11
0 26
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5523 0 0
2
5.90137e-315 0
0
13 Logic Switch~
5 51 336 0 10 11
0 27 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3330 0 0
2
5.90137e-315 0
0
13 Logic Switch~
5 49 196 0 1 11
0 28
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3465 0 0
2
5.90137e-315 0
0
13 Logic Switch~
5 50 170 0 1 11
0 29
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8396 0 0
2
5.90137e-315 0
0
13 Logic Switch~
5 50 145 0 1 11
0 30
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3685 0 0
2
5.90137e-315 0
0
13 Logic Switch~
5 51 116 0 1 11
0 31
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7849 0 0
2
5.90137e-315 0
0
13 Logic Switch~
5 53 87 0 10 11
0 32 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6343 0 0
2
5.90137e-315 0
0
7 Ground~
168 439 135 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7376 0 0
2
45537.4 0
0
7 Ground~
168 395 432 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9156 0 0
2
5.90137e-315 0
0
9 2-In AND~
219 1050 417 0 3 22
0 9 10 13
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
5776 0 0
2
5.90137e-315 0
0
6 74LS85
106 732 544 0 14 29
0 3 4 5 6 2 2 2 33 2
34 2 16 15 14
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U7
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
7207 0 0
2
5.90137e-315 5.34643e-315
0
6 74LS85
106 737 671 0 14 29
0 2 2 7 8 2 2 35 2 16
15 14 11 12 36
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U6
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
4459 0 0
2
5.90137e-315 5.32571e-315
0
7 Ground~
168 851 540 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3760 0 0
2
5.90137e-315 5.30499e-315
0
7 Ground~
168 639 835 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
754 0 0
2
5.90137e-315 5.26354e-315
0
8 2-In OR~
219 875 692 0 3 22
0 11 12 10
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
9767 0 0
2
5.90137e-315 0
0
8 2-In OR~
219 867 236 0 3 22
0 18 17 9
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
7978 0 0
2
5.90137e-315 0
0
7 Ground~
168 634 368 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3142 0 0
2
5.90137e-315 0
0
7 Ground~
168 846 73 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3284 0 0
2
5.90137e-315 0
0
6 74LS85
106 732 204 0 14 29
0 2 2 7 8 2 2 2 2 21
20 19 37 18 17
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U4
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
659 0 0
2
5.90137e-315 0
0
6 74LS85
106 727 77 0 14 29
0 3 4 5 6 38 39 2 40 2
41 2 21 20 19
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U3
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
3800 0 0
2
5.90137e-315 0
0
14 Logic Display~
6 1134 399 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6792 0 0
2
5.90137e-315 0
0
12 Hex Display~
7 449 77 0 16 19
10 8 7 2 2 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3701 0 0
2
5.90137e-315 0
0
12 Hex Display~
7 521 77 0 18 19
10 6 5 4 3 0 0 0 0 0
0 1 1 0 1 1 0 1 2
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
6316 0 0
2
5.90137e-315 0
0
7 74LS283
152 448 328 0 14 29
0 2 2 2 28 2 2 2 22 23
42 43 7 8 2
0
0 0 4848 0
7 74LS283
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 512 1 0 0 0
1 U
8734 0 0
2
5.90137e-315 0
0
7 74LS283
152 338 167 0 14 29
0 29 30 31 32 24 25 26 27 2
3 4 5 6 23
0
0 0 4848 0
7 74LS283
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 0 1 0 0 0
1 U
7988 0 0
2
5.90137e-315 0
0
72
4 0 2 0 0 4096 0 25 0 0 2 2
440 101
439 101
1 3 2 0 0 4112 0 11 25 0 0 4
439 129
439 100
446 100
446 101
1 0 2 0 0 0 0 12 0 0 4 2
395 426
395 427
0 0 2 0 0 0 0 0 0 0 54 2
395 432
395 427
0 1 3 0 0 8192 0 0 23 17 0 3
596 140
596 50
695 50
0 2 4 0 0 8192 0 0 23 18 0 3
585 150
585 59
695 59
0 3 5 0 0 8192 0 0 23 19 0 3
574 160
574 68
695 68
0 4 6 0 0 8192 0 0 23 20 0 3
565 169
565 77
695 77
6 0 2 0 0 4096 0 27 0 0 54 2
416 337
302 337
5 0 2 0 0 0 0 27 0 0 54 2
416 328
302 328
3 0 2 0 0 0 0 27 0 0 54 2
416 310
302 310
2 0 2 0 0 0 0 27 0 0 54 4
416 301
307 301
307 302
302 302
1 0 2 0 0 0 0 27 0 0 54 2
416 292
302 292
5 0 2 0 0 0 0 14 0 0 15 3
700 553
640 553
640 562
6 0 2 0 0 0 0 14 0 0 32 3
700 562
640 562
640 571
8 0 2 0 0 0 0 15 0 0 32 2
705 707
639 707
0 1 3 0 0 8320 0 0 14 57 0 4
512 140
597 140
597 517
700 517
0 2 4 0 0 8320 0 0 14 58 0 4
518 150
586 150
586 526
700 526
0 3 5 0 0 8320 0 0 14 59 0 4
524 160
575 160
575 535
700 535
0 4 6 0 0 8320 0 0 14 60 0 4
530 169
565 169
565 544
700 544
6 0 2 0 0 0 0 15 0 0 32 2
705 689
639 689
5 0 2 0 0 0 0 15 0 0 32 2
705 680
639 680
0 3 7 0 0 8320 0 0 15 55 0 4
490 337
548 337
548 662
705 662
0 4 8 0 0 8320 0 0 15 56 0 4
483 346
530 346
530 671
705 671
3 1 9 0 0 8320 0 19 13 0 0 4
900 236
1018 236
1018 408
1026 408
3 2 10 0 0 8320 0 18 13 0 0 4
908 692
1018 692
1018 426
1026 426
12 1 11 0 0 4224 0 15 18 0 0 4
769 689
854 689
854 683
862 683
13 2 12 0 0 4224 0 15 18 0 0 4
769 698
854 698
854 701
862 701
3 1 13 0 0 4224 0 13 24 0 0 2
1071 417
1134 417
1 0 2 0 0 0 0 15 0 0 32 2
705 644
639 644
2 0 2 0 0 0 0 15 0 0 32 2
705 653
639 653
7 1 2 0 0 8320 0 14 17 0 0 3
700 571
639 571
639 829
11 1 2 0 0 0 0 14 16 0 0 5
764 535
838 535
838 526
851 526
851 534
9 1 2 0 0 0 0 14 16 0 0 3
764 517
851 517
851 534
14 11 14 0 0 8320 0 14 15 0 0 4
764 580
793 580
793 662
769 662
13 10 15 0 0 8320 0 14 15 0 0 4
764 571
782 571
782 653
769 653
12 9 16 0 0 8320 0 14 15 0 0 4
764 562
773 562
773 644
769 644
5 0 2 0 0 0 0 22 0 0 46 2
700 213
634 213
6 0 2 0 0 0 0 22 0 0 46 4
700 222
639 222
639 223
634 223
7 0 2 0 0 0 0 22 0 0 46 2
700 231
634 231
1 0 2 0 0 0 0 22 0 0 46 2
700 177
634 177
2 0 2 0 0 0 0 22 0 0 46 2
700 186
634 186
14 2 17 0 0 4224 0 22 19 0 0 4
764 240
846 240
846 245
854 245
13 1 18 0 0 4224 0 22 19 0 0 4
764 231
846 231
846 227
854 227
8 0 2 0 0 0 0 22 0 0 46 2
700 240
634 240
7 1 2 0 0 0 0 23 20 0 0 3
695 104
634 104
634 362
11 1 2 0 0 0 0 23 21 0 0 5
759 68
833 68
833 59
846 59
846 67
9 1 2 0 0 0 0 23 21 0 0 3
759 50
846 50
846 67
14 11 19 0 0 8320 0 23 22 0 0 4
759 113
796 113
796 195
764 195
13 10 20 0 0 8320 0 23 22 0 0 4
759 104
785 104
785 186
764 186
12 9 21 0 0 8320 0 23 22 0 0 4
759 95
773 95
773 177
764 177
0 3 7 0 0 0 0 0 22 55 0 2
490 195
700 195
0 4 8 0 0 0 0 0 22 56 0 2
485 204
700 204
14 9 2 0 0 0 0 27 28 0 0 6
480 373
484 373
484 427
302 427
302 212
306 212
12 2 7 0 0 0 0 27 25 0 0 5
480 337
490 337
490 114
452 114
452 101
13 1 8 0 0 0 0 27 25 0 0 5
480 346
485 346
485 109
458 109
458 101
10 4 3 0 0 0 0 28 26 0 0 3
370 158
512 158
512 101
11 3 4 0 0 0 0 28 26 0 0 3
370 167
518 167
518 101
12 2 5 0 0 0 0 28 26 0 0 3
370 176
524 176
524 101
13 1 6 0 0 0 0 28 26 0 0 3
370 185
530 185
530 101
7 0 2 0 0 0 0 27 0 0 54 2
416 346
302 346
1 8 22 0 0 12416 0 1 27 0 0 4
62 443
192 443
192 355
416 355
14 9 23 0 0 8320 0 28 27 0 0 4
370 212
389 212
389 373
416 373
1 5 24 0 0 8320 0 2 28 0 0 4
61 420
141 420
141 167
306 167
1 6 25 0 0 8320 0 3 28 0 0 4
63 390
162 390
162 176
306 176
1 7 26 0 0 8320 0 4 28 0 0 4
64 361
175 361
175 185
306 185
1 8 27 0 0 8320 0 5 28 0 0 4
63 336
189 336
189 194
306 194
1 4 28 0 0 8320 0 6 27 0 0 5
61 196
61 212
271 212
271 319
416 319
1 1 29 0 0 12416 0 7 28 0 0 5
62 170
106 170
106 130
306 130
306 131
1 2 30 0 0 8320 0 8 28 0 0 3
62 145
62 140
306 140
1 3 31 0 0 12416 0 9 28 0 0 4
63 116
91 116
91 149
306 149
1 4 32 0 0 12416 0 10 28 0 0 4
65 87
74 87
74 158
306 158
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
