CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1358 699
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
76546066 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 399 35 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7901 0 0
2
5.90138e-315 0
0
13 Logic Switch~
5 466 36 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-8 -27 6 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4571 0 0
2
5.90138e-315 0
0
7 Ground~
168 568 567 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7796 0 0
2
5.90138e-315 0
0
7 74LS153
119 460 428 0 14 29
0 13 14 15 16 7 8 9 10 11
12 2 2 6 5
0
0 0 4848 0
7 74LS153
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 0 1 0 0 0
1 U
3907 0 0
2
5.90138e-315 0
0
7 74LS153
119 457 202 0 14 29
0 21 22 23 24 7 8 17 18 19
20 2 2 3 4
0
0 0 4848 0
7 74LS153
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 0 1 0 0 0
1 U
4389 0 0
2
5.90138e-315 0
0
8 Hex Key~
166 320 45 0 11 12
0 21 17 13 9 0 0 0 0 0
9 57
0
0 0 4656 0
0
4 KPD4
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
7762 0 0
2
5.90138e-315 0
0
8 Hex Key~
166 258 44 0 11 12
0 22 18 14 10 0 0 0 0 0
8 56
0
0 0 4656 0
0
4 KPD3
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
6723 0 0
2
5.90138e-315 0
0
8 Hex Key~
166 186 43 0 11 12
0 23 19 15 11 0 0 0 0 0
6 54
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
6871 0 0
2
5.90138e-315 0
0
12 Hex Display~
7 628 274 0 18 19
10 3 4 6 5 0 0 0 0 0
0 1 0 1 1 1 1 1 6
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4198 0 0
2
5.90138e-315 0
0
8 Hex Key~
166 109 44 0 11 12
0 24 20 16 12 0 0 0 0 0
9 57
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
970 0 0
2
5.90138e-315 0
0
28
11 0 2 0 0 4096 0 4 0 0 4 2
498 392
568 392
12 0 2 0 0 0 0 4 0 0 4 2
498 473
568 473
12 0 2 0 0 0 0 5 0 0 4 4
495 247
563 247
563 248
568 248
11 1 2 0 0 8320 0 5 3 0 0 3
495 166
568 166
568 561
13 1 3 0 0 8320 0 5 9 0 0 5
489 184
529 184
529 306
637 306
637 298
14 2 4 0 0 12416 0 5 9 0 0 5
489 229
514 229
514 321
631 321
631 298
14 4 5 0 0 8320 0 4 9 0 0 4
492 455
620 455
620 298
619 298
13 3 6 0 0 4224 0 4 9 0 0 3
492 410
625 410
625 298
0 5 7 0 0 8320 0 0 4 10 0 4
403 199
404 199
404 428
428 428
1 5 7 0 0 0 0 1 5 0 0 4
411 35
403 35
403 202
425 202
0 6 8 0 0 4224 0 0 4 12 0 3
376 210
376 437
428 437
1 6 8 0 0 0 0 2 5 0 0 5
478 36
478 110
376 110
376 211
425 211
4 7 9 0 0 4224 0 6 4 0 0 3
311 69
311 446
428 446
4 8 10 0 0 4224 0 7 4 0 0 3
249 68
249 455
428 455
4 9 11 0 0 4224 0 8 4 0 0 3
177 67
177 464
428 464
4 10 12 0 0 4224 0 10 4 0 0 3
100 68
100 473
428 473
3 1 13 0 0 4224 0 6 4 0 0 3
317 69
317 392
428 392
3 2 14 0 0 4224 0 7 4 0 0 3
255 68
255 401
428 401
3 3 15 0 0 4224 0 8 4 0 0 3
183 67
183 410
428 410
3 4 16 0 0 4224 0 10 4 0 0 3
106 68
106 419
428 419
2 7 17 0 0 4224 0 6 5 0 0 3
323 69
323 220
425 220
2 8 18 0 0 8320 0 7 5 0 0 3
261 68
261 229
425 229
2 9 19 0 0 8320 0 8 5 0 0 3
189 67
189 238
425 238
2 10 20 0 0 8320 0 10 5 0 0 3
112 68
112 247
425 247
1 1 21 0 0 4224 0 6 5 0 0 3
329 69
329 166
425 166
1 2 22 0 0 8320 0 7 5 0 0 3
267 68
267 175
425 175
1 3 23 0 0 8320 0 8 5 0 0 3
195 67
195 184
425 184
1 4 24 0 0 8320 0 10 5 0 0 3
118 68
118 193
425 193
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
