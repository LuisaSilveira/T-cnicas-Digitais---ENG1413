CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1358 699
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
76546066 0
0
6 Title:
5 Name:
0
0
0
15
13 Logic Switch~
5 92 384 0 1 11
0 10
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3409 0 0
2
45530.3 0
0
13 Logic Switch~
5 91 329 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3951 0 0
2
45530.3 1
0
13 Logic Switch~
5 90 266 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8885 0 0
2
45530.3 2
0
13 Logic Switch~
5 91 194 0 1 11
0 8
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3780 0 0
2
45530.3 3
0
13 Logic Switch~
5 91 129 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9265 0 0
2
45530.3 4
0
9 Inverter~
13 208 333 0 2 22
0 6 2
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 4 0
1 U
9442 0 0
2
45530.3 5
0
9 Inverter~
13 208 266 0 2 22
0 7 3
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 4 0
1 U
9424 0 0
2
45530.3 6
0
9 Inverter~
13 206 202 0 2 22
0 8 4
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
9968 0 0
2
45530.3 7
0
9 Inverter~
13 204 129 0 2 22
0 9 5
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
9281 0 0
2
45530.3 8
0
14 Logic Display~
6 826 293 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8464 0 0
2
45530.3 9
0
8 2-In OR~
219 701 328 0 3 22
0 13 12 11
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 18
65 0 0 0 4 1 5 0
1 U
7168 0 0
2
45530.3 10
0
8 2-In OR~
219 519 258 0 3 22
0 15 14 13
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 18
65 0 0 0 4 2 5 0
1 U
3171 0 0
2
45530.3 11
0
9 4-In AND~
219 343 430 0 5 22
0 5 4 3 2 12
0
0 0 608 0
6 74LS21
-21 -28 21 -20
3 U2A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 2 0
1 U
4139 0 0
2
45530.3 12
0
9 3-In AND~
219 343 329 0 4 22
0 3 2 10 14
0
0 0 608 0
6 74LS11
-21 -28 21 -20
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 1 0
1 U
6435 0 0
2
45530.3 13
0
9 3-In AND~
219 342 202 0 4 22
0 9 8 7 15
0
0 0 608 0
6 74LS11
-21 -28 21 -20
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 1 0
1 U
5283 0 0
2
45530.3 14
0
19
0 4 2 0 0 4224 0 0 13 5 0 3
236 329
236 444
319 444
0 3 3 0 0 4224 0 0 13 7 0 3
262 266
262 435
319 435
2 2 4 0 0 8320 0 8 13 0 0 4
227 202
283 202
283 426
319 426
2 1 5 0 0 8320 0 9 13 0 0 4
225 129
297 129
297 417
319 417
2 2 2 0 0 0 0 6 14 0 0 3
229 333
229 329
319 329
1 1 6 0 0 8320 0 2 6 0 0 3
103 329
103 333
193 333
2 1 3 0 0 0 0 7 14 0 0 4
229 266
311 266
311 320
319 320
0 3 7 0 0 8320 0 0 15 12 0 5
141 266
141 237
317 237
317 211
318 211
0 2 8 0 0 12416 0 0 15 13 0 6
143 202
144 202
144 226
310 226
310 202
318 202
0 1 9 0 0 8320 0 0 15 14 0 5
141 129
141 157
310 157
310 193
318 193
1 3 10 0 0 4224 0 1 14 0 0 4
104 384
311 384
311 338
319 338
1 1 7 0 0 0 0 3 7 0 0 2
102 266
193 266
1 1 8 0 0 0 0 4 8 0 0 3
103 194
103 202
191 202
1 1 9 0 0 0 0 5 9 0 0 2
103 129
189 129
3 1 11 0 0 4224 0 11 10 0 0 3
734 328
826 328
826 311
5 2 12 0 0 4224 0 13 11 0 0 4
364 430
680 430
680 337
688 337
3 1 13 0 0 4224 0 12 11 0 0 4
552 258
680 258
680 319
688 319
4 2 14 0 0 4224 0 14 12 0 0 4
364 329
498 329
498 267
506 267
1 4 15 0 0 4224 0 12 15 0 0 4
506 249
371 249
371 202
363 202
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
52 367 81 391
62 375 70 391
1 E
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
55 313 84 337
65 321 73 337
1 D
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
53 247 82 271
63 255 71 271
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
53 179 82 203
63 187 71 203
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
53 114 82 138
63 122 71 138
1 A
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
