CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 200 30 90 10
176 80 1358 699
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
76546066 0
0
6 Title:
5 Name:
0
0
0
42
13 Logic Switch~
5 56 825 0 10 11
0 41 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V14
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
469 0 0
2
45544.4 13
0
13 Logic Switch~
5 110 824 0 1 11
0 45
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V12
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4529 0 0
2
45544.4 12
0
13 Logic Switch~
5 157 824 0 1 11
0 44
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V11
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
88 0 0
2
45544.4 11
0
13 Logic Switch~
5 209 824 0 10 11
0 43 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3894 0 0
2
45544.4 10
0
13 Logic Switch~
5 261 823 0 10 11
0 42 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6890 0 0
2
45544.4 9
0
13 Logic Switch~
5 275 285 0 10 11
0 53 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3257 0 0
2
5.90138e-315 0
0
13 Logic Switch~
5 223 286 0 10 11
0 54 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6612 0 0
2
5.90138e-315 0
0
13 Logic Switch~
5 171 286 0 1 11
0 55
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3556 0 0
2
5.90138e-315 0
0
13 Logic Switch~
5 124 286 0 1 11
0 56
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9143 0 0
2
5.90138e-315 0
0
13 Logic Switch~
5 70 287 0 10 11
0 52 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8186 0 0
2
5.90138e-315 0
0
7 Ground~
168 874 954 0 1 3
0 2
0
0 0 53360 0
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3754 0 0
2
45544.5 0
0
12 Hex Display~
7 1866 616 0 18 19
10 9 8 7 6 0 0 0 0 0
0 1 1 1 1 1 1 1 8
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
8708 0 0
2
45544.4 0
0
12 Hex Display~
7 1775 618 0 18 19
10 13 11 10 12 0 0 0 0 0
0 1 1 1 1 0 0 1 3
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3338 0 0
2
45544.4 0
0
7 74LS283
152 1612 904 0 14 29
0 2 2 14 15 2 2 2 2 17
12 10 11 13 62
0
0 0 4848 0
7 74LS283
-24 -60 25 -52
3 U12
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 512 0 0 0 0
1 U
5546 0 0
2
45544.4 0
0
7 Ground~
168 1452 1059 0 1 3
0 2
0
0 0 53360 0
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3295 0 0
2
45544.4 0
0
7 74LS283
152 1528 723 0 14 29
0 21 20 19 18 2 22 22 2 16
6 7 8 9 17
0
0 0 4848 0
7 74LS283
-24 -60 25 -52
3 U11
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 0 0 0 0 0
1 U
4923 0 0
2
45544.4 0
0
7 Ground~
168 1206 917 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3248 0 0
2
45544.4 0
0
2 +V
167 1167 680 0 1 3
0 23
0
0 0 54256 0
2 5V
-7 -22 7 -14
3 V15
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3139 0 0
2
45544.4 0
0
7 Ground~
168 1327 556 0 1 3
0 2
0
0 0 53360 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3285 0 0
2
45544.4 3
0
2 +V
167 1296 620 0 1 3
0 24
0
0 0 54256 270
2 5V
-7 -15 7 -7
3 V16
-11 -25 10 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
336 0 0
2
45544.4 2
0
6 74LS85
106 1257 804 0 14 29
0 2 2 2 3 2 2 2 2 27
26 25 63 64 22
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
3 U14
-10 -62 11 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 0 0 0 0
1 U
6582 0 0
2
45544.4 1
0
6 74LS85
106 1254 637 0 14 29
0 21 20 19 18 23 2 2 23 2
24 2 27 26 25
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
3 U13
-10 -62 11 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 0 0 0 0 0
1 U
3546 0 0
2
45544.4 0
0
7 74LS283
152 974 791 0 14 29
0 2 2 28 29 2 2 30 31 3
65 66 14 15 16
0
0 0 4848 0
7 74LS283
-24 -60 25 -52
3 U10
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 512 0 0 0 0
1 U
893 0 0
2
45544.4 0
0
7 74LS283
152 973 610 0 14 29
0 36 37 38 39 32 33 34 35 2
21 20 19 18 3
0
0 0 4848 0
7 74LS283
-24 -60 25 -52
2 U9
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 0 0 0 0 0
1 U
8998 0 0
2
45544.4 0
0
6 74LS85
106 487 908 0 14 29
0 45 44 43 42 4 2 2 4 2
47 2 50 49 48
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U8
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 0 0 0 0 0
1 U
5979 0 0
2
45544.4 8
0
6 74LS85
106 490 1075 0 14 29
0 2 2 2 41 2 2 2 2 50
49 48 67 68 46
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U7
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 0 0 0 0
1 U
3835 0 0
2
45544.4 7
0
2 +V
167 386 1015 0 1 3
0 4
0
0 0 54256 0
2 5V
-5 -23 9 -15
2 V8
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
750 0 0
2
45544.4 6
0
7 Ground~
168 418 1171 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
849 0 0
2
45544.4 5
0
7 74LS283
152 654 914 0 14 29
0 45 44 43 42 2 46 46 2 2
32 33 34 35 40
0
0 0 4848 0
7 74LS283
-24 -60 25 -52
2 U4
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 0 0 0 0 0
1 U
4693 0 0
2
45544.4 4
0
7 74LS283
152 653 1078 0 14 29
0 2 2 2 41 2 2 2 2 40
69 70 30 31 71
0
0 0 4848 0
7 74LS283
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 512 0 0 0 0
1 U
4775 0 0
2
45544.4 3
0
2 +V
167 529 891 0 1 3
0 47
0
0 0 54256 270
2 5V
-7 -15 7 -7
2 V7
-8 -25 6 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9572 0 0
2
45544.4 2
0
7 Ground~
168 560 827 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3761 0 0
2
45544.4 1
0
7 Ground~
168 603 1195 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6765 0 0
2
45544.4 0
0
7 Ground~
168 617 657 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7938 0 0
2
45544.4 0
0
7 Ground~
168 574 289 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
55 0 0
2
45544.4 0
0
2 +V
167 543 353 0 1 3
0 58
0
0 0 54256 270
2 5V
-7 -15 7 -7
3 V13
-11 -25 10 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5610 0 0
2
45544.4 0
0
7 74LS283
152 667 540 0 14 29
0 2 2 2 52 2 2 2 2 51
72 73 28 29 74
0
0 0 4848 0
7 74LS283
-24 -60 25 -52
2 U6
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 512 0 0 0 0
1 U
3322 0 0
2
45544.4 0
0
7 74LS283
152 668 376 0 14 29
0 56 55 54 53 2 57 57 2 2
36 37 38 39 51
0
0 0 4848 0
7 74LS283
-24 -60 25 -52
2 U5
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 0 0 0 0 0
1 U
5914 0 0
2
45544.4 0
0
7 Ground~
168 432 633 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8748 0 0
2
45544.4 0
0
2 +V
167 400 477 0 1 3
0 5
0
0 0 54256 90
2 5V
-7 -15 7 -7
2 V1
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5830 0 0
2
45544.4 0
0
6 74LS85
106 504 537 0 14 29
0 2 2 2 52 2 2 2 2 61
60 59 75 76 57
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U3
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 0 0 0 0
1 U
9153 0 0
2
45544.4 0
0
6 74LS85
106 501 370 0 14 29
0 56 55 54 53 5 2 2 5 2
58 2 61 60 59
0
0 0 5104 0
6 74LS85
-21 -52 21 -44
2 U1
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 0 0 0 0 0
1 U
9220 0 0
2
45544.4 0
0
146
6 0 2 0 0 4096 0 23 0 0 5 2
942 800
874 800
5 0 2 0 0 0 0 23 0 0 5 4
942 791
879 791
879 792
874 792
2 0 2 0 0 0 0 23 0 0 5 2
942 764
874 764
1 0 2 0 0 0 0 23 0 0 5 2
942 755
874 755
9 1 2 0 0 8192 0 24 11 0 0 3
941 655
874 655
874 948
0 9 3 0 0 8320 0 0 23 7 0 4
1010 707
904 707
904 836
942 836
14 4 3 0 0 0 0 24 21 0 0 6
1005 655
1010 655
1010 707
1116 707
1116 804
1225 804
8 0 4 0 0 4096 0 25 0 0 105 2
455 944
386 944
8 0 5 0 0 4224 0 42 0 0 141 2
469 406
400 406
3 0 2 0 0 0 0 26 0 0 104 2
458 1066
418 1066
2 0 2 0 0 0 0 26 0 0 104 2
458 1057
418 1057
1 0 2 0 0 0 0 26 0 0 104 2
458 1048
418 1048
3 0 2 0 0 0 0 41 0 0 140 4
472 528
437 528
437 529
432 529
2 0 2 0 0 0 0 41 0 0 140 2
472 519
432 519
1 0 2 0 0 0 0 41 0 0 140 2
472 510
432 510
10 4 6 0 0 4224 0 16 12 0 0 3
1560 714
1857 714
1857 640
11 3 7 0 0 4224 0 16 12 0 0 3
1560 723
1863 723
1863 640
12 2 8 0 0 4224 0 16 12 0 0 3
1560 732
1869 732
1869 640
13 1 9 0 0 4224 0 16 12 0 0 3
1560 741
1875 741
1875 640
11 3 10 0 0 8320 0 14 13 0 0 3
1644 904
1772 904
1772 642
12 2 11 0 0 8320 0 14 13 0 0 3
1644 913
1778 913
1778 642
10 4 12 0 0 8320 0 14 13 0 0 3
1644 895
1766 895
1766 642
13 1 13 0 0 8320 0 14 13 0 0 3
1644 922
1784 922
1784 642
2 0 2 0 0 0 0 14 0 0 25 3
1580 877
1537 877
1537 868
1 0 2 0 0 0 0 14 0 0 35 2
1580 868
1452 868
12 3 14 0 0 12416 0 23 14 0 0 6
1006 800
1080 800
1080 885
1498 885
1498 886
1580 886
13 4 15 0 0 12416 0 23 14 0 0 4
1006 809
1063 809
1063 895
1580 895
14 9 16 0 0 12416 0 23 16 0 0 6
1006 836
1023 836
1023 861
1470 861
1470 768
1496 768
8 0 2 0 0 0 0 14 0 0 35 4
1580 931
1457 931
1457 932
1452 932
7 0 2 0 0 0 0 14 0 0 35 2
1580 922
1452 922
5 0 2 0 0 0 0 14 0 0 35 2
1580 904
1452 904
6 0 2 0 0 0 0 14 0 0 35 4
1580 913
1457 913
1457 914
1452 914
14 9 17 0 0 8320 0 16 14 0 0 4
1560 768
1572 768
1572 949
1580 949
8 0 2 0 0 0 0 16 0 0 35 2
1496 750
1452 750
5 1 2 0 0 8320 0 16 15 0 0 3
1496 723
1452 723
1452 1053
0 4 18 0 0 8320 0 0 16 53 0 5
1122 637
1122 533
1451 533
1451 714
1496 714
0 3 19 0 0 8320 0 0 16 54 0 5
1109 628
1109 521
1462 521
1462 705
1496 705
0 2 20 0 0 8320 0 0 16 55 0 5
1088 619
1088 509
1475 509
1475 696
1496 696
0 1 21 0 0 8320 0 0 16 56 0 5
1072 610
1072 499
1488 499
1488 687
1496 687
0 7 22 0 0 4224 0 0 16 41 0 2
1372 741
1496 741
14 6 22 0 0 0 0 21 16 0 0 4
1289 840
1372 840
1372 732
1496 732
8 0 2 0 0 0 0 21 0 0 50 2
1225 840
1206 840
7 0 2 0 0 0 0 21 0 0 50 2
1225 831
1206 831
6 0 2 0 0 0 0 21 0 0 50 2
1225 822
1206 822
5 0 2 0 0 0 0 21 0 0 50 2
1225 813
1206 813
3 0 2 0 0 0 0 21 0 0 50 2
1225 795
1206 795
2 0 2 0 0 0 0 21 0 0 50 2
1225 786
1206 786
1 0 2 0 0 0 0 21 0 0 50 4
1225 777
1211 777
1211 778
1206 778
7 0 2 0 0 0 0 22 0 0 50 2
1222 664
1206 664
6 1 2 0 0 0 0 22 17 0 0 3
1222 655
1206 655
1206 911
8 0 23 0 0 8320 0 22 0 0 52 4
1222 673
1222 711
1167 711
1167 696
5 1 23 0 0 128 0 22 18 0 0 5
1222 646
1192 646
1192 696
1167 696
1167 689
13 4 18 0 0 0 0 24 22 0 0 3
1005 628
1005 637
1222 637
12 3 19 0 0 0 0 24 22 0 0 4
1005 619
1015 619
1015 628
1222 628
11 2 20 0 0 0 0 24 22 0 0 4
1005 610
1025 610
1025 619
1222 619
10 1 21 0 0 0 0 24 22 0 0 4
1005 601
1033 601
1033 610
1222 610
11 0 2 0 0 0 0 22 0 0 58 3
1286 628
1313 628
1313 610
9 1 2 0 0 0 0 22 19 0 0 5
1286 610
1313 610
1313 542
1327 542
1327 550
1 10 24 0 0 4224 0 20 22 0 0 2
1284 619
1286 619
14 11 25 0 0 8320 0 22 21 0 0 4
1286 673
1307 673
1307 795
1289 795
13 10 26 0 0 8320 0 22 21 0 0 4
1286 664
1302 664
1302 786
1289 786
12 9 27 0 0 8320 0 22 21 0 0 4
1286 655
1297 655
1297 777
1289 777
12 3 28 0 0 8320 0 37 23 0 0 4
699 549
724 549
724 773
942 773
13 4 29 0 0 12416 0 37 23 0 0 4
699 558
714 558
714 782
942 782
12 7 30 0 0 8320 0 30 23 0 0 4
685 1087
929 1087
929 809
942 809
13 8 31 0 0 8320 0 30 23 0 0 4
685 1096
934 1096
934 818
942 818
10 5 32 0 0 8320 0 29 24 0 0 4
686 905
776 905
776 610
941 610
11 6 33 0 0 8320 0 29 24 0 0 4
686 914
783 914
783 619
941 619
12 7 34 0 0 8320 0 29 24 0 0 4
686 923
797 923
797 628
941 628
13 8 35 0 0 8320 0 29 24 0 0 4
686 932
811 932
811 637
941 637
10 1 36 0 0 8320 0 38 24 0 0 4
700 367
803 367
803 574
941 574
11 2 37 0 0 8320 0 38 24 0 0 4
700 376
792 376
792 583
941 583
12 3 38 0 0 8320 0 38 24 0 0 4
700 385
781 385
781 592
941 592
13 4 39 0 0 8320 0 38 24 0 0 4
700 394
773 394
773 601
941 601
14 9 40 0 0 16512 0 29 30 0 0 6
686 959
706 959
706 981
613 981
613 1123
621 1123
0 4 41 0 0 8192 0 0 30 106 0 5
334 1075
334 1138
583 1138
583 1069
621 1069
3 0 2 0 0 0 0 30 0 0 86 2
621 1060
603 1060
2 0 2 0 0 0 0 30 0 0 86 2
621 1051
603 1051
1 0 2 0 0 0 0 30 0 0 86 2
621 1042
603 1042
5 0 2 0 0 0 0 30 0 0 86 2
621 1078
603 1078
6 0 2 0 0 0 0 30 0 0 86 2
621 1087
603 1087
7 0 2 0 0 0 0 30 0 0 86 2
621 1096
603 1096
8 0 2 0 0 0 0 30 0 0 86 2
621 1105
603 1105
9 0 2 0 0 0 0 29 0 0 86 2
622 959
603 959
8 0 2 0 0 0 0 29 0 0 86 2
622 941
603 941
5 1 2 0 0 0 0 29 33 0 0 3
622 914
603 914
603 1189
0 4 42 0 0 8320 0 0 29 110 0 5
345 908
345 788
589 788
589 905
622 905
0 3 43 0 0 8320 0 0 29 109 0 5
359 899
359 776
598 776
598 896
622 896
0 2 44 0 0 8192 0 0 29 108 0 5
370 890
370 762
607 762
607 887
622 887
0 1 45 0 0 8192 0 0 29 107 0 5
383 881
383 751
614 751
614 878
622 878
0 7 46 0 0 4096 0 0 29 92 0 4
573 935
614 935
614 932
622 932
14 6 46 0 0 8320 0 26 29 0 0 4
522 1111
573 1111
573 923
622 923
11 0 2 0 0 0 0 25 0 0 94 3
519 899
546 899
546 881
9 1 2 0 0 0 0 25 32 0 0 5
519 881
546 881
546 813
560 813
560 821
1 10 47 0 0 4224 0 31 25 0 0 2
517 890
519 890
14 11 48 0 0 8320 0 25 26 0 0 4
519 944
540 944
540 1066
522 1066
13 10 49 0 0 8320 0 25 26 0 0 4
519 935
535 935
535 1057
522 1057
12 9 50 0 0 8320 0 25 26 0 0 4
519 926
530 926
530 1048
522 1048
7 0 2 0 0 0 0 25 0 0 104 2
455 935
418 935
8 0 2 0 0 0 0 26 0 0 104 2
458 1111
418 1111
7 0 2 0 0 0 0 26 0 0 104 2
458 1102
418 1102
6 0 2 0 0 0 0 26 0 0 104 2
458 1093
418 1093
5 0 2 0 0 0 0 26 0 0 104 2
458 1084
418 1084
6 1 2 0 0 0 0 25 28 0 0 4
455 926
455 925
418 925
418 1165
5 1 4 0 0 8320 0 25 27 0 0 3
455 917
386 917
386 1024
1 4 41 0 0 12416 0 1 26 0 0 4
68 825
85 825
85 1075
458 1075
1 1 45 0 0 12416 0 2 25 0 0 4
122 824
132 824
132 881
455 881
1 2 44 0 0 12416 0 3 25 0 0 4
169 824
184 824
184 890
455 890
1 3 43 0 0 0 0 4 25 0 0 4
221 824
237 824
237 899
455 899
1 4 42 0 0 0 0 5 25 0 0 4
273 823
281 823
281 908
455 908
14 9 51 0 0 16512 0 38 37 0 0 6
700 421
720 421
720 443
627 443
627 585
635 585
0 4 52 0 0 8192 0 0 37 142 0 5
348 537
348 600
597 600
597 531
635 531
3 0 2 0 0 0 0 37 0 0 122 2
635 522
617 522
2 0 2 0 0 0 0 37 0 0 122 2
635 513
617 513
1 0 2 0 0 0 0 37 0 0 122 2
635 504
617 504
5 0 2 0 0 0 0 37 0 0 122 2
635 540
617 540
6 0 2 0 0 0 0 37 0 0 122 2
635 549
617 549
7 0 2 0 0 0 0 37 0 0 122 2
635 558
617 558
8 0 2 0 0 0 0 37 0 0 122 2
635 567
617 567
9 0 2 0 0 0 0 38 0 0 122 2
636 421
617 421
8 0 2 0 0 0 0 38 0 0 122 2
636 403
617 403
5 1 2 0 0 0 0 38 34 0 0 3
636 376
617 376
617 651
0 4 53 0 0 8320 0 0 38 146 0 5
359 370
359 250
603 250
603 367
636 367
0 3 54 0 0 8320 0 0 38 145 0 5
373 361
373 238
612 238
612 358
636 358
0 2 55 0 0 8192 0 0 38 144 0 5
384 352
384 224
621 224
621 349
636 349
0 1 56 0 0 8192 0 0 38 143 0 5
397 343
397 213
628 213
628 340
636 340
0 7 57 0 0 4096 0 0 38 128 0 4
587 395
628 395
628 394
636 394
14 6 57 0 0 8320 0 41 38 0 0 4
536 573
587 573
587 385
636 385
11 0 2 0 0 0 0 42 0 0 130 3
533 361
560 361
560 343
9 1 2 0 0 0 0 42 35 0 0 5
533 343
560 343
560 275
574 275
574 283
1 10 58 0 0 4224 0 36 42 0 0 2
531 352
533 352
14 11 59 0 0 8320 0 42 41 0 0 4
533 406
554 406
554 528
536 528
13 10 60 0 0 8320 0 42 41 0 0 4
533 397
549 397
549 519
536 519
12 9 61 0 0 8320 0 42 41 0 0 4
533 388
544 388
544 510
536 510
7 0 2 0 0 0 0 42 0 0 140 2
469 397
432 397
8 0 2 0 0 0 0 41 0 0 140 2
472 573
432 573
7 0 2 0 0 0 0 41 0 0 140 2
472 564
432 564
6 0 2 0 0 0 0 41 0 0 140 2
472 555
432 555
5 0 2 0 0 0 0 41 0 0 140 2
472 546
432 546
6 1 2 0 0 0 0 42 39 0 0 4
469 388
469 389
432 389
432 627
5 1 5 0 0 144 0 42 40 0 0 6
469 379
400 379
400 411
419 411
419 475
411 475
1 4 52 0 0 12416 0 10 41 0 0 4
82 287
99 287
99 537
472 537
1 1 56 0 0 12416 0 9 42 0 0 4
136 286
146 286
146 343
469 343
1 2 55 0 0 12416 0 8 42 0 0 4
183 286
198 286
198 352
469 352
1 3 54 0 0 0 0 7 42 0 0 4
235 286
251 286
251 361
469 361
1 4 53 0 0 0 0 6 42 0 0 4
287 285
295 285
295 370
469 370
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
